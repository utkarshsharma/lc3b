// alu.vh - ALU header file

`ifndef _alu_vh_
`define _alu_vh_

// ALU operations
`define alu_add 2'b00 // a + b
`define alu_and 2'b01 // a & b
`define alu_xor 2'b10 // a ^ b
`define alu_a   2'b11 // a

`endif //_alu_vh_
