`ifndef _pc_vh_
`define _pc_vh_

`define PCMUX_INC  2'b00 // PC + 2
`define PCMUX_BUS  2'b01 // value from bus
`define PCMUX_ADDR 2'b10 // output from address adder

`define PC_RST 16'b0 // PC reset value

`endif //_pc_vh_
